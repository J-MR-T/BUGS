module _4zmbitz_DEC (clk, rst, Enable, Input_1, Input_2, Input_3, Input_4, Output_1, Output_2, Output_3, Output_4, Output_5, Output_6, Output_7, Output_8, Output_9, Output_10, Output_11, Output_12, Output_13, Output_14, Output_15, Output_16);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Enable;
  input  wire [0:0] Input_1;
  input  wire [0:0] Input_2;
  input  wire [0:0] Input_3;
  input  wire [0:0] Input_4;
  output  wire [0:0] Output_1;
  output  wire [0:0] Output_2;
  output  wire [0:0] Output_3;
  output  wire [0:0] Output_4;
  output  wire [0:0] Output_5;
  output  wire [0:0] Output_6;
  output  wire [0:0] Output_7;
  output  wire [0:0] Output_8;
  output  wire [0:0] Output_9;
  output  wire [0:0] Output_10;
  output  wire [0:0] Output_11;
  output  wire [0:0] Output_12;
  output  wire [0:0] Output_13;
  output  wire [0:0] Output_14;
  output  wire [0:0] Output_15;
  output  wire [0:0] Output_16;

  TC_Decoder3 # (.UUID(64'd3557036857616701976 ^ UUID)) Decoder3_0 (.dis(wire_3), .sel0(wire_11), .sel1(wire_1), .sel2(wire_4), .out0(wire_22), .out1(wire_13), .out2(wire_7), .out3(wire_0), .out4(wire_19), .out5(wire_10), .out6(wire_9), .out7(wire_25));
  TC_Decoder3 # (.UUID(64'd3820282478237721292 ^ UUID)) Decoder3_1 (.dis(wire_21), .sel0(wire_11), .sel1(wire_1), .sel2(wire_4), .out0(wire_24), .out1(wire_18), .out2(wire_23), .out3(wire_20), .out4(wire_8), .out5(wire_5), .out6(wire_16), .out7(wire_14));
  TC_Not # (.UUID(64'd4201052158732111988 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_6), .out(wire_12));
  TC_And # (.UUID(64'd4454436996045823864 ^ UUID), .BIT_WIDTH(64'd1)) And_3 (.in0(wire_2), .in1(wire_12), .out(wire_17));
  TC_And # (.UUID(64'd4393166029961138605 ^ UUID), .BIT_WIDTH(64'd1)) And_4 (.in0(wire_2), .in1(wire_6), .out(wire_15));
  TC_Not # (.UUID(64'd3447179360407859019 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_15), .out(wire_3));
  TC_Not # (.UUID(64'd89992856383661183 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_17), .out(wire_21));

  wire [0:0] wire_0;
  assign Output_2 = wire_0;
  wire [0:0] wire_1;
  assign wire_1 = Input_2;
  wire [0:0] wire_2;
  assign wire_2 = Enable;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  assign wire_4 = Input_3;
  wire [0:0] wire_5;
  assign Output_12 = wire_5;
  wire [0:0] wire_6;
  assign wire_6 = Input_4;
  wire [0:0] wire_7;
  assign Output_1 = wire_7;
  wire [0:0] wire_8;
  assign Output_11 = wire_8;
  wire [0:0] wire_9;
  assign Output_5 = wire_9;
  wire [0:0] wire_10;
  assign Output_8 = wire_10;
  wire [0:0] wire_11;
  assign wire_11 = Input_1;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  assign Output_4 = wire_13;
  wire [0:0] wire_14;
  assign Output_10 = wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  assign Output_9 = wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  assign Output_16 = wire_18;
  wire [0:0] wire_19;
  assign Output_7 = wire_19;
  wire [0:0] wire_20;
  assign Output_14 = wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  assign Output_3 = wire_22;
  wire [0:0] wire_23;
  assign Output_13 = wire_23;
  wire [0:0] wire_24;
  assign Output_15 = wire_24;
  wire [0:0] wire_25;
  assign Output_6 = wire_25;

endmodule
