module BUGS (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Switch # (.UUID(64'd2889093244921319772 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_0 (.en(wire_31), .in(wire_113), .out(wire_5_3));
  TC_Switch # (.UUID(64'd86943380849751926 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_1 (.en(wire_122), .in(wire_106), .out(wire_5_2));
  TC_Switch # (.UUID(64'd4014842671027375889 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_2 (.en(wire_129), .in(wire_33), .out(wire_5_1));
  TC_Switch # (.UUID(64'd61774588077662089 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_118), .in(wire_16), .out(wire_5_0));
  TC_Switch # (.UUID(64'd2259330822597661583 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_123), .in(wire_113), .out(wire_15_0));
  TC_Switch # (.UUID(64'd45211650065772438 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_120), .in(wire_106), .out(wire_15_1));
  TC_Switch # (.UUID(64'd636641294393885960 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_127), .in(wire_33), .out(wire_15_2));
  TC_Switch # (.UUID(64'd1187325688266991947 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_78), .in(wire_16), .out(wire_15_3));
  TC_Splitter16 # (.UUID(64'd2786955280030538084 ^ UUID)) Splitter16_8 (.in(wire_94[15:0]), .out0(wire_99), .out1(wire_73));
  TC_Splitter8 # (.UUID(64'd1512558103295404783 ^ UUID)) Splitter8_9 (.in(wire_99), .out0(wire_57), .out1(wire_46), .out2(wire_102), .out3(wire_104), .out4(wire_67), .out5(wire_25), .out6(wire_77), .out7(wire_49));
  TC_Splitter8 # (.UUID(64'd2739075887445410243 ^ UUID)) Splitter8_10 (.in(wire_73), .out0(), .out1(), .out2(), .out3(), .out4(wire_72), .out5(wire_11), .out6(wire_91), .out7(wire_112));
  TC_Program # (.UUID(64'd1962896349348883544 ^ UUID), .WORD_WIDTH(64'd16), .DEFAULT_FILE_NAME("Program_1B3D9BD471D9EC58.w16.bin"), .ARG_SIG("Program_1B3D9BD471D9EC58=%s")) Program_11 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_0 }), .out0(wire_94), .out1(), .out2(), .out3());
  TC_Maker8 # (.UUID(64'd1811210392590479892 ^ UUID)) Maker8_12 (.in0(wire_67), .in1(wire_25), .in2(wire_77), .in3(wire_49), .in4(wire_49), .in5(wire_49), .in6(wire_49), .in7(wire_49), .out(wire_28));
  TC_Switch # (.UUID(64'd59861540961676004 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_3), .in(wire_135), .out(wire_4_3));
  TC_Decoder3 # (.UUID(64'd1091720397448825704 ^ UUID)) Decoder3_14 (.dis(1'd0), .sel0(wire_11), .sel1(wire_91), .sel2(wire_112), .out0(wire_32), .out1(wire_3), .out2(wire_74), .out3(wire_13), .out4(wire_21), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd284066621739992948 ^ UUID)) Splitter8_15 (.in(wire_73), .out0(wire_64), .out1(wire_27), .out2(wire_96), .out3(wire_125), .out4(), .out5(), .out6(), .out7());
  TC_And3 # (.UUID(64'd2349936586489369383 ^ UUID), .BIT_WIDTH(64'd1)) And3_16 (.in0(wire_64), .in1(wire_27), .in2(wire_95), .out(wire_58));
  TC_Not # (.UUID(64'd1862029186245978007 ^ UUID), .BIT_WIDTH(64'd1)) Not_17 (.in(wire_125), .out(wire_19));
  TC_Not # (.UUID(64'd2886023162162490038 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_96), .out(wire_95));
  TC_Not # (.UUID(64'd4547963649571443974 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_131), .out(wire_128));
  TC_Add # (.UUID(64'd2219056279148372749 ^ UUID), .BIT_WIDTH(64'd8)) Add8_20 (.in0({{7{1'b0}}, wire_14 }), .in1(wire_0), .ci(1'd0), .out(wire_52), .co());
  TC_Constant # (.UUID(64'd284927449043062334 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_21 (.out(wire_14));
  TC_Mux # (.UUID(64'd1490074330709799775 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_22 (.sel(wire_26), .in0(wire_52), .in1(wire_5), .out(wire_40));
  TC_And # (.UUID(64'd4571478384267617773 ^ UUID), .BIT_WIDTH(64'd1)) And_23 (.in0(wire_58), .in1(wire_19), .out(wire_131));
  TC_Mux # (.UUID(64'd4390152381466029418 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_24 (.sel(wire_133), .in0(wire_28), .in1(wire_15), .out(wire_44));
  TC_Not # (.UUID(64'd739297898705157967 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_72), .out(wire_133));
  TC_Splitter8 # (.UUID(64'd2346719092904309270 ^ UUID)) Splitter8_26 (.in(wire_73), .out0(wire_65), .out1(wire_37), .out2(wire_86), .out3(wire_134), .out4(), .out5(), .out6(), .out7());
  TC_And # (.UUID(64'd2778597424498181009 ^ UUID), .BIT_WIDTH(64'd1)) And_27 (.in0(wire_71), .in1(wire_74), .out(wire_26));
  TC_Maker8 # (.UUID(64'd272098822319972058 ^ UUID)) Maker8_28 (.in0(wire_130), .in1(wire_69), .in2(wire_132), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_48));
  TC_Splitter8 # (.UUID(64'd3610426648490400219 ^ UUID)) Splitter8_29 (.in(wire_48), .out0(wire_8), .out1(wire_17), .out2(wire_63), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3482878620302494581 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_30 (.en(wire_107), .in(wire_17), .out(wire_23_9));
  TC_Switch # (.UUID(64'd3634901032405140120 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_31 (.en(wire_43), .in(wire_116), .out(wire_23_8));
  TC_Not # (.UUID(64'd1546046292452294576 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_17), .out(wire_116));
  TC_Switch # (.UUID(64'd2992728460288496718 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_33 (.en(wire_90), .in(wire_92), .out(wire_23_6));
  TC_And # (.UUID(64'd967663677127503883 ^ UUID), .BIT_WIDTH(64'd1)) And_34 (.in0(wire_59), .in1(wire_22), .out(wire_92));
  TC_Not # (.UUID(64'd330724126800016971 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_63), .out(wire_10));
  TC_Not # (.UUID(64'd4153118730818407170 ^ UUID), .BIT_WIDTH(64'd1)) Not_36 (.in(wire_17), .out(wire_59));
  TC_Not # (.UUID(64'd248193864262529728 ^ UUID), .BIT_WIDTH(64'd1)) Not_37 (.in(wire_8), .out(wire_22));
  TC_Switch # (.UUID(64'd1256931279237961986 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_38 (.en(wire_45), .in(wire_8), .out(wire_23_4));
  TC_Switch # (.UUID(64'd1565021323724993591 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_39 (.en(wire_42), .in(wire_22), .out(wire_23_2));
  TC_Switch # (.UUID(64'd1741380941796187096 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_40 (.en(wire_51), .in(wire_105), .out(wire_23_0));
  TC_Or # (.UUID(64'd638524781242385127 ^ UUID), .BIT_WIDTH(64'd1)) Or_41 (.in0(wire_17), .in1(wire_8), .out(wire_105));
  TC_Switch # (.UUID(64'd259266863711477162 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_42 (.en(wire_66), .in(wire_63), .out(wire_23_1));
  TC_Switch # (.UUID(64'd2305268859645322721 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_43 (.en(wire_47), .in(wire_126), .out(wire_23_3));
  TC_And # (.UUID(64'd3718192804095311357 ^ UUID), .BIT_WIDTH(64'd1)) And_44 (.in0(wire_59), .in1(wire_10), .out(wire_126));
  TC_Switch # (.UUID(64'd3258303036381579932 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_45 (.en(wire_60), .in(wire_119), .out(wire_23_5));
  TC_Or # (.UUID(64'd39189119703468738 ^ UUID), .BIT_WIDTH(64'd1)) Or_46 (.in0(wire_17), .in1(wire_63), .out(wire_119));
  TC_Switch # (.UUID(64'd3829403973650022461 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_47 (.en(wire_89), .in(wire_10), .out(wire_23_7));
  TC_Or # (.UUID(64'd2278039841302013877 ^ UUID), .BIT_WIDTH(64'd1)) Or_48 (.in0(wire_79), .in1(wire_117), .out(wire_62));
  TC_And # (.UUID(64'd2848714878388336043 ^ UUID), .BIT_WIDTH(64'd1)) And_49 (.in0(wire_128), .in1(wire_3), .out(wire_108));
  TC_Or3 # (.UUID(64'd2418308136627262819 ^ UUID), .BIT_WIDTH(64'd1)) Or3_50 (.in0(wire_23), .in1(wire_79), .in2(wire_97), .out(wire_71));
  TC_Splitter8 # (.UUID(64'd3227541871505226795 ^ UUID)) Splitter8_51 (.in(wire_93), .out0(), .out1(), .out2(wire_36), .out3(wire_35), .out4(wire_7), .out5(wire_136), .out6(wire_83), .out7(wire_109));
  TC_Splitter8 # (.UUID(64'd4082558212404249919 ^ UUID)) Splitter8_52 (.in(wire_68), .out0(wire_110), .out1(wire_24), .out2(wire_12), .out3(wire_103), .out4(), .out5(), .out6(), .out7());
  TC_Splitter16 # (.UUID(64'd3854874253491533690 ^ UUID)) Splitter16_53 (.in(wire_94[15:0]), .out0(wire_93), .out1(wire_68));
  TC_Maker8 # (.UUID(64'd4135035395817306410 ^ UUID)) Maker8_54 (.in0(wire_7), .in1(wire_136), .in2(wire_83), .in3(wire_109), .in4(wire_110), .in5(wire_24), .in6(wire_12), .in7(wire_103), .out(wire_84));
  TC_And # (.UUID(64'd2870407041976778370 ^ UUID), .BIT_WIDTH(64'd1)) And_55 (.in0(wire_3), .in1(wire_108), .out(wire_56));
  TC_Switch # (.UUID(64'd2373468547285715425 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_56 (.en(wire_79), .in(wire_52), .out(wire_4_1));
  TC_Switch # (.UUID(64'd4280956778265416790 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_57 (.en(wire_13), .in(wire_84), .out(wire_4_2));
  TC_Ram # (.UUID(64'd3749859122203513419 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd65536)) Ram_58 (.clk(clk), .rst(rst), .load(wire_29), .save(wire_53), .address({{16{1'b0}}, wire_82 }), .in0({{56{1'b0}}, wire_9 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_20), .out1(), .out2(), .out3());
  TC_Maker16 # (.UUID(64'd2412269050531193143 ^ UUID)) Maker16_59 (.in0(wire_5), .in1(wire_15), .out(wire_61));
  TC_Decoder1 # (.UUID(64'd2739246431798704612 ^ UUID)) Decoder1_60 (.sel(wire_72), .out0(wire_100), .out1(wire_41));
  TC_Switch # (.UUID(64'd659273495617936174 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_61 (.en(wire_29), .in(wire_20[7:0]), .out(wire_4_0));
  TC_Or3 # (.UUID(64'd4081227845994135766 ^ UUID), .BIT_WIDTH(64'd1)) Or3_62 (.in0(wire_13), .in1(wire_29), .in2(wire_56), .out(wire_85));
  TC_Not # (.UUID(64'd737816774998180178 ^ UUID), .BIT_WIDTH(64'd1)) Not_63 (.in(wire_29), .out(wire_87));
  TC_Switch # (.UUID(64'd50166919081845044 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_64 (.en(wire_30), .in(wire_16), .out(wire_9_0));
  TC_Switch # (.UUID(64'd256379383749359748 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_65 (.en(wire_38), .in(wire_33), .out(wire_9_1));
  TC_Switch # (.UUID(64'd3361432240314569015 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_66 (.en(wire_98), .in(wire_106), .out(wire_9_3));
  TC_Switch # (.UUID(64'd2326822053092830863 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_67 (.en(wire_88), .in(wire_113), .out(wire_9_2));
  TC_Switch # (.UUID(64'd7233660929838003 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_68 (.en(wire_21), .in(wire_100), .out(wire_29));
  TC_Switch # (.UUID(64'd270113544502984811 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_69 (.en(wire_21), .in(wire_41), .out(wire_53));
  TC_Or # (.UUID(64'd3847373968220149442 ^ UUID), .BIT_WIDTH(64'd1)) Or_70 (.in0(wire_3), .in1(wire_21), .out(wire_75));
  TC_Or3 # (.UUID(64'd1164534403528806362 ^ UUID), .BIT_WIDTH(64'd1)) Or3_71 (.in0(wire_3), .in1(wire_21), .in2(wire_74), .out(wire_124));
  TC_Maker8 # (.UUID(64'd1108719941909561335 ^ UUID)) Maker8_72 (.in0(wire_55), .in1(wire_81), .in2(wire_65), .in3(wire_37), .in4(wire_86), .in5(wire_134), .in6(1'd0), .in7(1'd0), .out(wire_6));
  TC_Splitter8 # (.UUID(64'd4492080329498477228 ^ UUID)) Splitter8_73 (.in(wire_99), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(), .out6(wire_55), .out7(wire_81));
  TC_Add # (.UUID(64'd2078765471029358326 ^ UUID), .BIT_WIDTH(64'd16)) Add16_74 (.in0(wire_61), .in1(wire_80), .ci(1'd0), .out(wire_82), .co());
  TC_Splitter8 # (.UUID(64'd1560050035605001328 ^ UUID)) Splitter8_75 (.in(wire_6), .out0(wire_18), .out1(wire_39), .out2(wire_137), .out3(wire_114), .out4(wire_121), .out5(wire_1), .out6(), .out7());
  TC_Maker8 # (.UUID(64'd2888961188701163738 ^ UUID)) Maker8_76 (.in0(wire_18), .in1(wire_39), .in2(wire_137), .in3(wire_114), .in4(wire_121), .in5(wire_1), .in6(wire_1), .in7(wire_1), .out(wire_111));
  TC_Maker8 # (.UUID(64'd241675556150898430 ^ UUID)) Maker8_77 (.in0(wire_1), .in1(wire_1), .in2(wire_1), .in3(wire_1), .in4(wire_1), .in5(wire_1), .in6(wire_1), .in7(wire_1), .out(wire_101));
  TC_Maker16 # (.UUID(64'd2957865413649645104 ^ UUID)) Maker16_78 (.in0(wire_111), .in1(wire_101), .out(wire_80));
  WEz_Reg8 # (.UUID(64'd582847863739762236 ^ UUID)) WEz_Reg8_79 (.clk(clk), .rst(rst), .Input(wire_4), .Write_Enable(wire_34), .Output(wire_113));
  WEz_Reg8 # (.UUID(64'd2457469979817797657 ^ UUID)) WEz_Reg8_80 (.clk(clk), .rst(rst), .Input(wire_4), .Write_Enable(wire_76), .Output(wire_106));
  WEz_Reg8 # (.UUID(64'd1658420752031332203 ^ UUID)) WEz_Reg8_81 (.clk(clk), .rst(rst), .Input(wire_4), .Write_Enable(wire_54), .Output(wire_33));
  WEz_Reg8 # (.UUID(64'd1645122552538795091 ^ UUID)) WEz_Reg8_82 (.clk(clk), .rst(rst), .Input(wire_4), .Write_Enable(wire_62), .Output(wire_16));
  _2zmbitz_DEC # (.UUID(64'd2197142114939782149 ^ UUID)) _2zmbitz_DEC_83 (.clk(clk), .rst(rst), .Upper(wire_25), .Lower(wire_67), .Enable(wire_75), .\3 (wire_78), .\0 (wire_123), .\1 (wire_120), .\2 (wire_127));
  _2zmbitz_DEC # (.UUID(64'd1549555523845691351 ^ UUID)) _2zmbitz_DEC_84 (.clk(clk), .rst(rst), .Upper(wire_46), .Lower(wire_57), .Enable(wire_85), .\3 (wire_117), .\0 (wire_34), .\1 (wire_76), .\2 (wire_54));
  _2zmbitz_DEC # (.UUID(64'd2027745803572602827 ^ UUID)) _2zmbitz_DEC_85 (.clk(clk), .rst(rst), .Upper(wire_104), .Lower(wire_102), .Enable(wire_124), .\3 (wire_118), .\0 (wire_31), .\1 (wire_122), .\2 (wire_129));
  WEz_Reg8 # (.UUID(64'd1907960194756986957 ^ UUID)) WEz_Reg8_86 (.clk(clk), .rst(rst), .Input(wire_40), .Write_Enable(wire_14), .Output(wire_0));
  ALU2 # (.UUID(64'd3726698497104897986 ^ UUID)) ALU2_87 (.clk(clk), .rst(rst), .Input_1(wire_5), .Input_2(wire_44), .Instruction(wire_73), .\ALU? (wire_3), .CF(wire_130), .ZF(wire_69), .SF(wire_132), .Output(wire_135));
  _4zmbitz_DEC # (.UUID(64'd3551504769601007530 ^ UUID)) _4zmbitz_DEC_88 (.clk(clk), .rst(rst), .Enable(wire_74), .Input_1(wire_65), .Input_2(wire_37), .Input_3(wire_86), .Input_4(wire_134), .Output_1(wire_60), .Output_2(wire_89), .Output_3(wire_66), .Output_4(wire_47), .Output_5(wire_2), .Output_6(wire_50), .Output_7(wire_115), .Output_8(wire_70), .Output_9(wire_42), .Output_10(wire_51), .Output_11(wire_90), .Output_12(wire_45), .Output_13(wire_107), .Output_14(wire_43), .Output_15(wire_97), .Output_16(wire_79));
  _2zmbitz_DEC # (.UUID(64'd74734672557308173 ^ UUID)) _2zmbitz_DEC_89 (.clk(clk), .rst(rst), .Upper(wire_46), .Lower(wire_57), .Enable(wire_87), .\3 (wire_30), .\0 (wire_88), .\1 (wire_98), .\2 (wire_38));

  wire [7:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_4_0;
  wire [7:0] wire_4_1;
  wire [7:0] wire_4_2;
  wire [7:0] wire_4_3;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3;
  wire [7:0] wire_5;
  wire [7:0] wire_5_0;
  wire [7:0] wire_5_1;
  wire [7:0] wire_5_2;
  wire [7:0] wire_5_3;
  assign wire_5 = wire_5_0|wire_5_1|wire_5_2|wire_5_3;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_9_0;
  wire [7:0] wire_9_1;
  wire [7:0] wire_9_2;
  wire [7:0] wire_9_3;
  assign wire_9 = wire_9_0|wire_9_1|wire_9_2|wire_9_3;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_15_0;
  wire [7:0] wire_15_1;
  wire [7:0] wire_15_2;
  wire [7:0] wire_15_3;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2|wire_15_3;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [63:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_23_0;
  wire [0:0] wire_23_1;
  wire [0:0] wire_23_2;
  wire [0:0] wire_23_3;
  wire [0:0] wire_23_4;
  wire [0:0] wire_23_5;
  wire [0:0] wire_23_6;
  wire [0:0] wire_23_7;
  wire [0:0] wire_23_8;
  wire [0:0] wire_23_9;
  assign wire_23 = wire_23_0|wire_23_1|wire_23_2|wire_23_3|wire_23_4|wire_23_5|wire_23_6|wire_23_7|wire_23_8|wire_23_9;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [7:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [15:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [15:0] wire_80;
  wire [0:0] wire_81;
  wire [15:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [7:0] wire_93;
  wire [63:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [7:0] wire_99;
  wire [0:0] wire_100;
  wire [7:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [7:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [7:0] wire_111;
  wire [0:0] wire_112;
  wire [7:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [0:0] wire_126;
  wire [0:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [0:0] wire_131;
  wire [0:0] wire_132;
  wire [0:0] wire_133;
  wire [0:0] wire_134;
  wire [7:0] wire_135;
  wire [0:0] wire_136;
  wire [0:0] wire_137;

endmodule
